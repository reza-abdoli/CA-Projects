module instructionMemory(A,RD);
input [31:0] A;
output reg [31:0] RD;
reg [31:0] mem [64000:0];
initial begin
$readmemh("program.txt",mem);
end
always @ (*) begin
 	 RD = mem[A[31:2]];
end

endmodule

